module dLatch
  
endmodule


module dFlipflop
  
  
endmodule 
